** sch_path: /secondary/opt/pdk/lf11_xschem/lf11_pdk_xschem/test_mosLF_4_7.sch
**.subckt test_mosLF_4_7
V1 VG 0 0.3
V2 VD 0 0.5
V3 net2 0 1.2
V4 net3 0 0.7
V5 net1 0 0.95
xm1 net3 net1 net2 net2 pmos1v2hvt L=0.11e-6 W=1e-6 nf=1 abdrain='int((nf+1)/2) * W/nf * 0.30e-6' absource='int((nf+2)/2) * W/nf * 0.30e-6'
+ lsdrain='2*int((nf+1)/2) * (W/nf + 0.30e-6)' lssource='2*int((nf+2)/2) * (W/nf + 0.30e-6)' dta=0 nrd='0.30e-6 / W' nrs='0.30e-6 / W'
+ sa=0.36e-6 sb=0.36e-6 sd=0 mult=1 m=1
xm2 VD VG 0 0 nmos1v2hvt L=0.11e-6 W=1e-6 nf=1 abdrain='int((nf+1)/2) * W/nf * 0.30e-6' absource='int((nf+2)/2) * W/nf * 0.30e-6' lsdrain='2*int((nf+1)/2) * (W/nf + 0.30e-6)'
+ lssource='2*int((nf+2)/2) * (W/nf + 0.30e-6)' dta=0 nrd='0.30e-6 / W' nrs='0.30e-6 / W' sa=0.36e-6 sb=0.36e-6 sd=0 mult=1 m=1
**** begin user architecture code


.lib '../../../models/montecarlo_config.lib' mc_off
.lib '../../../models/lf11is.lib' 1v2hvt_tt

.option temp=27
.option savecurrents
.save all @n.xm1.nm1[gm] @n.xm1.nm1[ids] @n.xm2.nm1[gm] @n.xm2.nm1[ids]

.control
pre_osdi ../../../models/psp103.osdi
op
write test_mosLF_4_7.raw
.endc


**** end user architecture code
**.ends
.end
