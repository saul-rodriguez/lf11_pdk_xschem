** sch_path: /secondary/opt/pdk/lf11_xschem/lf11_pdk_xschem/test_cmimsLF.sch
**.subckt test_cmimsLF
XC1 net1 0 cmims w=33e-6 l=33e-6 m=1
V1 net1 0 1
**** begin user architecture code


.lib '../../../models/lf11is.lib' mim_typ
*Following lines necessary for DcOp
.option savecurrents
.save all
*
.control
*DcOp
op
write rc_filter.raw

.endc


**** end user architecture code
**.ends
.end
